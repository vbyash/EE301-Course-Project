magic
tech scmos
timestamp 1699134136
<< nwell >>
rect -126 142 372 189
rect -127 26 372 142
<< ntransistor >>
rect -31 -17 -27 -13
rect 140 -16 144 -14
rect 162 -16 262 -14
rect 296 -16 327 -14
rect 139 -58 144 -56
rect 191 -60 211 -56
rect 296 -60 327 -58
<< ptransistor >>
rect -103 81 49 83
rect 252 110 264 112
rect 105 81 172 83
rect 200 80 206 84
rect 237 58 277 60
<< ndiffusion >>
rect -31 -3 -27 1
rect -31 -13 -27 -8
rect 140 -14 144 -2
rect 162 -8 205 1
rect 216 -8 262 1
rect 162 -14 262 -8
rect 296 -3 310 1
rect 316 -3 327 1
rect 296 -14 327 -3
rect -31 -22 -27 -17
rect 140 -22 144 -16
rect 162 -23 262 -16
rect -31 -31 -27 -27
rect 162 -31 205 -23
rect 216 -31 262 -23
rect 296 -27 327 -16
rect 296 -31 310 -27
rect 316 -31 327 -27
rect 139 -46 144 -41
rect 139 -56 144 -51
rect 191 -48 199 -41
rect 204 -48 211 -41
rect 191 -56 211 -48
rect 296 -47 310 -42
rect 316 -47 327 -42
rect 139 -63 144 -58
rect 296 -58 327 -47
rect 139 -73 144 -68
rect 191 -66 211 -60
rect 191 -73 199 -66
rect 204 -73 211 -66
rect 296 -69 327 -60
rect 296 -74 310 -69
rect 316 -74 327 -69
<< pdiffusion >>
rect 252 124 264 131
rect -103 90 -40 124
rect -13 90 49 124
rect 105 98 129 122
rect 150 98 172 122
rect -103 83 49 90
rect 105 83 172 98
rect 200 114 206 122
rect 252 112 264 118
rect 200 84 206 106
rect 252 104 264 110
rect 252 91 264 98
rect -103 73 49 81
rect -103 40 -40 73
rect -13 40 49 73
rect 105 67 172 81
rect 105 40 129 67
rect 150 40 172 67
rect 200 55 206 80
rect 237 70 255 80
rect 262 70 277 80
rect 237 60 277 70
rect 200 40 206 47
rect 237 50 277 58
rect 237 40 255 50
rect 262 40 277 50
<< ndcontact >>
rect -31 -8 -27 -3
rect 140 -2 144 3
rect 205 -8 216 1
rect 310 -3 316 1
rect -31 -27 -27 -22
rect 140 -27 144 -22
rect 205 -31 216 -23
rect 310 -31 316 -27
rect 139 -51 144 -46
rect 199 -48 204 -41
rect 310 -47 316 -42
rect 139 -68 144 -63
rect 199 -73 204 -66
rect 310 -74 316 -69
<< pdcontact >>
rect -40 90 -13 124
rect 129 98 150 122
rect 200 106 206 114
rect 252 118 264 124
rect 252 98 264 104
rect -40 40 -13 73
rect 129 40 150 67
rect 255 70 262 80
rect 200 47 206 55
rect 255 40 262 50
<< psubstratepcontact >>
rect -23 -113 -18 -90
rect 146 -113 150 -90
rect 199 -113 204 -90
rect 310 -113 316 -90
<< nsubstratencontact >>
rect -40 156 -13 177
rect 129 156 150 177
rect 210 156 216 177
rect 243 156 249 177
<< polysilicon >>
rect -107 81 -103 83
rect 49 81 57 83
rect 66 81 75 83
rect 84 81 90 83
rect 235 110 252 112
rect 264 110 270 112
rect 276 110 282 112
rect 99 81 105 83
rect 172 81 188 83
rect 193 80 200 84
rect 206 80 214 84
rect 223 58 227 60
rect 233 58 237 60
rect 277 58 291 60
rect -46 -17 -43 -13
rect -37 -17 -31 -13
rect -27 -17 -12 -13
rect 119 -16 126 -14
rect 132 -16 140 -14
rect 144 -16 162 -14
rect 262 -16 296 -14
rect 327 -16 343 -14
rect 119 -58 139 -56
rect 144 -58 155 -56
rect 177 -60 181 -56
rect 186 -60 191 -56
rect 211 -60 225 -56
rect 281 -60 286 -58
rect 291 -60 296 -58
rect 327 -60 339 -58
<< polycontact >>
rect 57 81 66 92
rect 90 81 99 92
rect 270 110 276 114
rect 214 80 219 84
rect 227 58 233 62
rect -43 -17 -37 -13
rect 126 -16 132 -12
rect 155 -58 159 -54
rect 181 -60 186 -56
rect 286 -60 291 -56
<< metal1 >>
rect -90 156 -40 177
rect -13 156 129 177
rect 150 156 210 177
rect 216 156 243 177
rect 249 156 280 177
rect -40 124 -13 156
rect 129 122 150 156
rect 75 100 82 106
rect 57 94 99 100
rect 210 114 216 156
rect 243 124 249 156
rect 243 118 252 124
rect 270 118 316 123
rect 206 106 216 114
rect 270 114 276 118
rect 310 114 316 118
rect 310 109 325 114
rect 222 101 228 107
rect 57 92 66 94
rect 90 92 99 94
rect 214 93 233 101
rect 214 84 219 93
rect 227 72 233 93
rect 245 98 252 104
rect 245 87 250 98
rect 245 82 262 87
rect 210 67 233 72
rect 255 80 262 82
rect -40 26 -13 40
rect 210 55 216 67
rect 227 62 233 67
rect 206 47 216 55
rect 129 30 150 40
rect -25 10 -19 26
rect -43 4 -19 10
rect -43 -13 -37 4
rect -25 -3 -19 4
rect 146 3 150 30
rect 209 9 216 47
rect 255 39 262 40
rect 310 39 316 109
rect 255 33 316 39
rect -27 -5 -19 -3
rect 68 -5 74 1
rect 144 2 150 3
rect 144 -2 159 2
rect -27 -8 132 -5
rect -25 -9 132 -8
rect 126 -12 132 -9
rect -27 -27 -18 -22
rect 144 -27 150 -22
rect -23 -90 -18 -27
rect 146 -46 150 -27
rect 144 -51 150 -46
rect 155 -47 159 -2
rect 205 1 216 9
rect 310 1 316 33
rect 205 -35 216 -31
rect 199 -40 216 -35
rect 199 -41 204 -40
rect 155 -51 186 -47
rect 310 -42 316 -31
rect 155 -54 159 -51
rect 181 -55 291 -51
rect 181 -56 186 -55
rect 286 -56 291 -55
rect 144 -68 150 -63
rect 146 -90 150 -68
rect 199 -90 204 -73
rect 310 -90 316 -74
rect -59 -113 -23 -90
rect -18 -113 146 -90
rect 150 -113 199 -90
rect 204 -113 310 -90
rect 316 -113 349 -90
<< labels >>
rlabel metal1 75 106 82 106 1 V_biasp
rlabel metal1 68 1 74 1 1 V_bias3
rlabel metal1 222 107 228 107 1 V_bias2
rlabel metal1 325 109 325 114 1 V_bias1
rlabel metal1 171 -99 171 -99 1 gnd
rlabel metal1 175 168 175 168 1 vdd
<< end >>
